library verilog;
use verilog.vl_types.all;
entity tf_test is
end tf_test;
