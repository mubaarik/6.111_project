// File:   zbt_6111_sample.v
// Date:   26-Nov-05
// Author: I. Chuang <ichuang@mit.edu>
//
// Sample code for the MIT 6.111 labkit demonstrating use of the ZBT
// memories for video display.  Video input from the NTSC digitizer is
// displayed within an XGA 1024x768 window.  One ZBT memory (ram0) is used
// as the video frame buffer, with 8 bits used per pixel (black & white).
//
// Since the ZBT is read once for every four pixels, this frees up time for 
// data to be stored to the ZBT during other pixel times.  The NTSC decoder
// runs at 27 MHz, whereas the XGA runs at 65 MHz, so we synchronize
// signals between the two (see ntsc2zbt.v) and let the NTSC data be
// stored to ZBT memory whenever it is available, during cycles when
// pixel reads are not being performed.
//
// We use a very simple ZBT interface, which does not involve any clock
// generation or hiding of the pipelining.  See zbt_6111.v for more info.
//
// switch[7] selects between display of NTSC video and test bars
// switch[6] is used for testing the NTSC decoder
// switch[1] selects between test bar periods; these are stored to ZBT
//           during blanking periods
// switch[0] selects vertical test bars (hardwired; not stored in ZBT)
//
//
// Bug fix: Jonathan P. Mailoa <jpmailoa@mit.edu>
// Date   : 11-May-09
////
// Use ramclock module to deskew clocks;  GPH
// To change display from 1024*787 to 800*600, use clock_40mhz and change
// accordingly. Verilog ntsc2zbt.v will also need changes to change resolution.
//
// Date   : 10-Nov-11

///////////////////////////////////////////////////////////////////////////////
//
// 6.111 FPGA Labkit -- Template Toplevel Module
//
// For Labkit Revision 004
//
//
// Created: October 31, 2004, from revision 003 file
// Author: Nathan Ickes
//
///////////////////////////////////////////////////////////////////////////////
//
//
// CHANGES FOR BOARD REVISION 004
//
// 1) Added signals for logic analyzer pods 2-4.
// 2) Expanded "tv_in_ycrcb" to 20 bits.
// 3) Renamed "tv_out_data" to "tv_out_i2c_data" and "tv_out_sclk" to
//    "tv_out_i2c_clock".
// 4) Reversed disp_data_in and disp_data_out signals, so that "out" is an
//    output of the FPGA, and "in" is an input.
//
// CHANGES FOR BOARD REVISION 003
//
// 1) Combined flash chip enables into a single signal, flash_ce_b.
//
// CHANGES FOR BOARD REVISION 002
//
// 1) Added SRAM clock feedback path input and output
// 2) Renamed "mousedata" to "mouse_data"
// 3) Renamed some ZBT memory signals. Parity bits are now incorporated into 
//    the data bus, and the byte write enables have been combined into the
//    4-bit ram#_bwe_b bus.
// 4) Removed the "systemace_clock" net, since the SystemACE clock is now
//    hardwired on the PCB to the oscillator.
//
///////////////////////////////////////////////////////////////////////////////
//
// Complete change history (including bug fixes)
//
// 2011-Nov-10: Changed resolution to 1024 * 768.
//					 Added back ramclok to deskew RAM clock
//
// 2009-May-11: Fixed memory management bug by 8 clock cycle forecast. 
//              Changed resolution to  800 * 600.
//              Reduced clock speed to 40MHz.
//              Disconnected zbt_6111's ram_clk signal. 
//              Added ramclock to control RAM.
//              Added notes about ram1 default values.
//              Commented out clock_feedback_out assignment.
//              Removed delayN modules because ZBT's latency has no more effect.
//
// 2005-Sep-09: Added missing default assignments to "ac97_sdata_out",
//              "disp_data_out", "analyzer[2-3]_clock" and
//              "analyzer[2-3]_data".
//
// 2005-Jan-23: Reduced flash address bus to 24 bits, to match 128Mb devices
//              actually populated on the boards. (The boards support up to
//              256Mb devices, with 25 address lines.)
//
// 2004-Oct-31: Adapted to new revision 004 board.
//
// 2004-May-01: Changed "disp_data_in" to be an output, and gave it a default
//              value. (Previous versions of this file declared this port to
//              be an input.)
//
// 2004-Apr-29: Reduced SRAM address busses to 19 bits, to match 18Mb devices
//              actually populated on the boards. (The boards support up to
//              72Mb devices, with 21 address lines.)
//
// 2004-Apr-29: Change history started
//
///////////////////////////////////////////////////////////////////////////////

module zbt_6111_sample(beep, audio_reset_b, 
		       ac97_sdata_out, ac97_sdata_in, ac97_synch,
	       ac97_bit_clock,
	       
	       vga_out_red, vga_out_green, vga_out_blue, vga_out_sync_b,
	       vga_out_blank_b, vga_out_pixel_clock, vga_out_hsync,
	       vga_out_vsync,

	       tv_out_ycrcb, tv_out_reset_b, tv_out_clock, tv_out_i2c_clock,
	       tv_out_i2c_data, tv_out_pal_ntsc, tv_out_hsync_b,
	       tv_out_vsync_b, tv_out_blank_b, tv_out_subcar_reset,

	       tv_in_ycrcb, tv_in_data_valid, tv_in_line_clock1,
	       tv_in_line_clock2, tv_in_aef, tv_in_hff, tv_in_aff,
	       tv_in_i2c_clock, tv_in_i2c_data, tv_in_fifo_read,
	       tv_in_fifo_clock, tv_in_iso, tv_in_reset_b, tv_in_clock,

	       ram0_data, ram0_address, ram0_adv_ld, ram0_clk, ram0_cen_b,
	       ram0_ce_b, ram0_oe_b, ram0_we_b, ram0_bwe_b, 

	       ram1_data, ram1_address, ram1_adv_ld, ram1_clk, ram1_cen_b,
	       ram1_ce_b, ram1_oe_b, ram1_we_b, ram1_bwe_b,

	       clock_feedback_out, clock_feedback_in,

	       flash_data, flash_address, flash_ce_b, flash_oe_b, flash_we_b,
	       flash_reset_b, flash_sts, flash_byte_b,

	       rs232_txd, rs232_rxd, rs232_rts, rs232_cts,

	       mouse_clock, mouse_data, keyboard_clock, keyboard_data,

	       clock_27mhz, clock1, clock2,

	       disp_blank, disp_data_out, disp_clock, disp_rs, disp_ce_b,
	       disp_reset_b, disp_data_in,

	       button0, button1, button2, button3, button_enter, button_right,
	       button_left, button_down, button_up,

	       switch,

	       led,
	       
	       user1, user2, user3, user4,
	       
	       daughtercard,

	       systemace_data, systemace_address, systemace_ce_b,
	       systemace_we_b, systemace_oe_b, systemace_irq, systemace_mpbrdy,
	       
	       analyzer1_data, analyzer1_clock,
 	       analyzer2_data, analyzer2_clock,
 	       analyzer3_data, analyzer3_clock,
 	       analyzer4_data, analyzer4_clock);

   output beep, audio_reset_b, ac97_synch, ac97_sdata_out;
   input  ac97_bit_clock, ac97_sdata_in;
   
   output [7:0] vga_out_red, vga_out_green, vga_out_blue;
   output vga_out_sync_b, vga_out_blank_b, vga_out_pixel_clock,
	  vga_out_hsync, vga_out_vsync;

   output [9:0] tv_out_ycrcb;
   output tv_out_reset_b, tv_out_clock, tv_out_i2c_clock, tv_out_i2c_data,
	  tv_out_pal_ntsc, tv_out_hsync_b, tv_out_vsync_b, tv_out_blank_b,
	  tv_out_subcar_reset;
   
   input  [19:0] tv_in_ycrcb;
   input  tv_in_data_valid, tv_in_line_clock1, tv_in_line_clock2, tv_in_aef,
	  tv_in_hff, tv_in_aff;
   output tv_in_i2c_clock, tv_in_fifo_read, tv_in_fifo_clock, tv_in_iso,
	  tv_in_reset_b, tv_in_clock;
   inout  tv_in_i2c_data;
        
   inout  [35:0] ram0_data;
   output [18:0] ram0_address;
   output ram0_adv_ld, ram0_clk, ram0_cen_b, ram0_ce_b, ram0_oe_b, ram0_we_b;
   output [3:0] ram0_bwe_b;
   
   inout  [35:0] ram1_data;
   output [18:0] ram1_address;
   output ram1_adv_ld, ram1_clk, ram1_cen_b, ram1_ce_b, ram1_oe_b, ram1_we_b;
   output [3:0] ram1_bwe_b;

   input  clock_feedback_in;
   output clock_feedback_out;
   
   inout  [15:0] flash_data;
   output [24:0] flash_address;
   output flash_ce_b, flash_oe_b, flash_we_b, flash_reset_b, flash_byte_b;
   input  flash_sts;
   
   output rs232_txd, rs232_rts;
   input  rs232_rxd, rs232_cts;

   input  mouse_clock, mouse_data, keyboard_clock, keyboard_data;

   input  clock_27mhz, clock1, clock2;

   output disp_blank, disp_clock, disp_rs, disp_ce_b, disp_reset_b;  
   input  disp_data_in;
   output  disp_data_out;
   
   input  button0, button1, button2, button3, button_enter, button_right,
	  button_left, button_down, button_up;
   input  [7:0] switch;
   output [7:0] led;

   inout [31:0] user1, user2, user3, user4;
   
   inout [43:0] daughtercard;

   inout  [15:0] systemace_data;
   output [6:0]  systemace_address;
   output systemace_ce_b, systemace_we_b, systemace_oe_b;
   input  systemace_irq, systemace_mpbrdy;

   output [15:0] analyzer1_data, analyzer2_data, analyzer3_data, 
		 analyzer4_data;
   output analyzer1_clock, analyzer2_clock, analyzer3_clock, analyzer4_clock;

   ////////////////////////////////////////////////////////////////////////////
   //
   // I/O Assignments
   //
   ////////////////////////////////////////////////////////////////////////////
   
   // Audio Input and Output
   assign beep= 1'b0;
   assign audio_reset_b = 1'b0;
   assign ac97_synch = 1'b0;
   assign ac97_sdata_out = 1'b0;
/*
*/
   // ac97_sdata_in is an input

   // Video Output
   assign tv_out_ycrcb = 10'h0;
   assign tv_out_reset_b = 1'b0;
   assign tv_out_clock = 1'b0;
   assign tv_out_i2c_clock = 1'b0;
   assign tv_out_i2c_data = 1'b0;
   assign tv_out_pal_ntsc = 1'b0;
   assign tv_out_hsync_b = 1'b1;
   assign tv_out_vsync_b = 1'b1;
   assign tv_out_blank_b = 1'b1;
   assign tv_out_subcar_reset = 1'b0;
   
   // Video Input
   //assign tv_in_i2c_clock = 1'b0;
   assign tv_in_fifo_read = 1'b1;
   assign tv_in_fifo_clock = 1'b0;
   assign tv_in_iso = 1'b1;
   //assign tv_in_reset_b = 1'b0;
   assign tv_in_clock = clock_27mhz;//1'b0;
   //assign tv_in_i2c_data = 1'bZ;
   // tv_in_ycrcb, tv_in_data_valid, tv_in_line_clock1, tv_in_line_clock2, 
   // tv_in_aef, tv_in_hff, and tv_in_aff are inputs
   
   // SRAMs

/* change lines below to enable ZBT RAM bank0 */

/*
   assign ram0_data = 36'hZ;
   assign ram0_address = 19'h0;
   assign ram0_clk = 1'b0;
   assign ram0_we_b = 1'b1;
   assign ram0_cen_b = 1'b0;	// clock enable
*/

/* enable RAM pins */

   assign ram0_ce_b = 1'b0;
   assign ram0_oe_b = 1'b0;
   assign ram0_adv_ld = 1'b0;
   assign ram0_bwe_b = 4'h0; 

/**********/

   assign ram1_data = 36'hZ; 
   assign ram1_address = 19'h0;
   assign ram1_adv_ld = 1'b0;
   assign ram1_clk = 1'b0;
   
   //These values has to be set to 0 like ram0 if ram1 is used.
   assign ram1_cen_b = 1'b1;
   assign ram1_ce_b = 1'b1;
   assign ram1_oe_b = 1'b1;
   assign ram1_we_b = 1'b1;
   assign ram1_bwe_b = 4'hF;

   // clock_feedback_out will be assigned by ramclock
   // assign clock_feedback_out = 1'b0;  //2011-Nov-10
   // clock_feedback_in is an input
   
   // Flash ROM
   assign flash_data = 16'hZ;
   assign flash_address = 25'h0;
   assign flash_ce_b = 1'b1;
   assign flash_oe_b = 1'b1;
   assign flash_we_b = 1'b1;
   assign flash_reset_b = 1'b0;
   assign flash_byte_b = 1'b1;
   // flash_sts is an input

   // RS-232 Interface
   assign rs232_txd = 1'b1;
   assign rs232_rts = 1'b1;
   // rs232_rxd and rs232_cts are inputs

   // PS/2 Ports
   // mouse_clock, mouse_data, keyboard_clock, and keyboard_data are inputs

   // LED Displays
/*
   assign disp_blank = 1'b1;
   assign disp_clock = 1'b0;
   assign disp_rs = 1'b0;
   assign disp_ce_b = 1'b1;
   assign disp_reset_b = 1'b0;
   assign disp_data_out = 1'b0;
*/
   // disp_data_in is an input

   // Buttons, Switches, and Individual LEDs
   //lab3 assign led = 8'hFF;
   // button0, button1, button2, button3, button_enter, button_right,
   // button_left, button_down, button_up, and switches are inputs

   // User I/Os
   assign user1 = 32'hZ;
   assign user2 = 32'hZ;
   assign user3 = 32'hZ;
   assign user4 = 32'hZ;

   // Daughtercard Connectors
   assign daughtercard = 44'hZ;

   // SystemACE Microprocessor Port
   assign systemace_data = 16'hZ;
   assign systemace_address = 7'h0;
   assign systemace_ce_b = 1'b1;
   assign systemace_we_b = 1'b1;
   assign systemace_oe_b = 1'b1;
   // systemace_irq and systemace_mpbrdy are inputs

   // Logic Analyzer
   assign analyzer1_data = 16'h0;
   assign analyzer1_clock = 1'b1;
   assign analyzer2_data = 16'h0;
   assign analyzer2_clock = 1'b1;
   //assign analyzer3_data = 16'h0;
   //assign analyzer3_clock = 1'b1;
   assign analyzer4_data = 16'h0;
   assign analyzer4_clock = 1'b1;
		    
   ////////////////////////////////////////////////////////////////////////////
   // Demonstration of ZBT RAM as video memory

   // use FPGA's digital clock manager to produce a
   // 65MHz clock (actually 64.8MHz)
   wire clock_65mhz_unbuf,clock_65mhz;
   DCM vclk1(.CLKIN(clock_27mhz),.CLKFX(clock_65mhz_unbuf));
   // synthesis attribute CLKFX_DIVIDE of vclk1 is 10
   // synthesis attribute CLKFX_MULTIPLY of vclk1 is 24
   // synthesis attribute CLK_FEEDBACK of vclk1 is NONE
   // synthesis attribute CLKIN_PERIOD of vclk1 is 37
   BUFG vclk2(.O(clock_65mhz),.I(clock_65mhz_unbuf));

//   wire clk = clock_65mhz;  // gph 2011-Nov-10

/*
   ////////////////////////////////////////////////////////////////////////////
   // Demonstration of ZBT RAM as video memory
   // use FPGA's digital clock manager to produce a
   // 40MHz clock (actually 40.5MHz)
   wire clock_40mhz_unbuf,clock_40mhz;
   DCM vclk1(.CLKIN(clock_27mhz),.CLKFX(clock_40mhz_unbuf));
   // synthesis attribute CLKFX_DIVIDE of vclk1 is 2
   // synthesis attribute CLKFX_MULTIPLY of vclk1 is 3
   // synthesis attribute CLK_FEEDBACK of vclk1 is NONE
   // synthesis attribute CLKIN_PERIOD of vclk1 is 37
   BUFG vclk2(.O(clock_40mhz),.I(clock_40mhz_unbuf));
//   wire clk = clock_40mhz;
*/

	wire locked;

	//assign clock_feedback_out = 0; // gph 2011-Nov-10
   
   ramclock rc(.ref_clock(clock_65mhz), .fpga_clock(clk),
					.ram0_clock(ram0_clk), 
					//.ram1_clock(ram1_clk),   //uncomment if ram1 is used
					.clock_feedback_in(clock_feedback_in),
					.clock_feedback_out(clock_feedback_out), .locked(locked));

   
   // power-on reset generation
   wire power_on_reset;    // remain high for first 16 clocks
   SRL16 reset_sr (.D(1'b0), .CLK(clk), .Q(power_on_reset),
		   .A0(1'b1), .A1(1'b1), .A2(1'b1), .A3(1'b1));
   defparam reset_sr.INIT = 16'hFFFF;

   // ENTER button is user reset
   wire reset,user_reset, trigger, clear;
   debounce db1(power_on_reset, clk, ~button_left, user_reset);
	debounce db2(power_on_reset, clk, ~user3[1], clear);
	debounce db3(power_on_reset, clk, user3[0], trigger);
   assign reset = user_reset | power_on_reset;
   
	
   // display module for debugging

   reg [63:0] dispdata;
   display_16hex hexdisp1(reset, clk, dispdata,
			  disp_blank, disp_clock, disp_rs, disp_ce_b,
			  disp_reset_b, disp_data_out);

   // generate basic XVGA video signals
   wire [10:0] hcount;
   wire [9:0]  vcount;
   wire hsync,vsync,blank;
   xvga xvga1(clk,hcount,vcount,hsync,vsync,blank);
   
	wire in_frame;
   assign in_frame = (hcount > 34) & (hcount < 744)
                   & (vcount > 78) & (vcount < 564);
   // wire up to ZBT ram

   wire [35:0] vram_write_data;
   wire [35:0] vram_read_data;
   wire [18:0] vram_addr;
   wire        vram_we;

   wire ram0_clk_not_used;
   zbt_6111 zbt1(clk, 1'b1, vram_we, vram_addr,
		   vram_write_data, vram_read_data,
		   ram0_clk_not_used,   //to get good timing, don't connect ram_clk to zbt_6111
		   ram0_we_b, ram0_address, ram0_data, ram0_cen_b);

   // generate pixel value from reading ZBT memory
   wire [17:0] 	vr_pixel;
   wire [18:0] 	vram_addr1;
   wire [10:0] center_x;
	wire [9:0] center_y;
	wire [31:0] whiteCount, sumX, sumY;
	wire divided, reseted, white;
   vram_display vd1(reset,clk,hcount,vcount,vr_pixel, center_x, center_y,whiteCount, sumX, sumY,reseted, divided,white,
		    vram_addr1,vram_read_data);

   // ADV7185 NTSC decoder interface code
   // adv7185 initialization module
   adv7185init adv7185(.reset(reset), .clock_27mhz(clock_27mhz), 
		       .source(1'b0), .tv_in_reset_b(tv_in_reset_b), 
		       .tv_in_i2c_clock(tv_in_i2c_clock), 
		       .tv_in_i2c_data(tv_in_i2c_data));

   wire [29:0] ycrcb;	// video data (luminance, chrominance)
   wire [2:0] fvh;	// sync for field, vertical, horizontal
   wire       dv;	// data valid
   
   ntsc_decode decode (.clk(tv_in_line_clock1), .reset(reset),
		       .tv_in_ycrcb(tv_in_ycrcb[19:10]), 
		       .ycrcb(ycrcb), .f(fvh[2]),
		       .v(fvh[1]), .h(fvh[0]), .data_valid(dv));

   reg [2:0] xfvh [1:0];
	reg xdv [1:0];
	
	always @(posedge clk) begin 
		{xfvh[1], xfvh[0]}={xfvh[0], fvh};
		{xdv[1],xdv[0]}={xdv[0], dv};
	end
   // convert ycrcb to RGB
   wire [7:0] R, G, B;
   wire [9:0] Y, Cr, Cb;
   assign Y = ycrcb[29:20];
   assign Cr = ycrcb[19:10];
   assign Cb = ycrcb[9:0];
   YCrCb2RGB rgb_conv ( .R(R), .G(G), .B(B), 
                        .clk(tv_in_line_clock1), .rst(0), 
                        .Y(Y), .Cr(Cr), .Cb(Cb) );
   //////HSV conversion here
	wire [7:0] _h,_s,_v, black_white;
	rgb2hsv hsv(.clock(clk), .reset(0), .r(R), .g(G), .b(B), .h(_h), ._s(_s), .v(_v));
	///////////////
	/////thresholding colors 
	///////////////
	wire [7:0] r_black_white, b_black_white, g_black_white, o_black_white; 
	//green
	hsv_thresh #(.h_high_thresh(150), .s_high_thresh(230), .v_high_thresh(255),.h_low_thresh(70), .s_low_thresh(80), .v_low_thresh(200))
	thresh (.clock(clk),.red(0), .reset(0), .H(_h), .S(_s), .V(_v), .color(g_black_white));
	//red
	hsv_thresh #(.h_high_thresh(255), .s_high_thresh(230), .v_high_thresh(255),.h_low_thresh(246), .s_low_thresh(80), .v_low_thresh(200))
	thresh1 (.clock(clk),.red(1), .reset(0), .H(_h), .S(_s), .V(_v), .color(r_black_white));
	//orange 
	hsv_thresh #(.h_high_thresh(35), .s_high_thresh(230), .v_high_thresh(255),.h_low_thresh(15), .s_low_thresh(80), .v_low_thresh(200))
	thresh2 (.clock(clk),.red(0), .reset(0), .H(_h), .S(_s), .V(_v), .color(o_black_white));
	//blue 
	hsv_thresh #(.h_high_thresh(170), .s_high_thresh(230), .v_high_thresh(255),.h_low_thresh(140), .s_low_thresh(80), .v_low_thresh(200))
	thresh3 (.clock(clk),.red(0), .reset(0), .H(_h), .S(_s), .V(_v), .color(b_black_white));
	////erosion
	//wire [7:0] erode = b_black_white+g_black_white+r_black_white+o_black_white;
	wire [7:0] dialated;
	//erosion e(.clock(clk),.reset(reset),.hcount(hcount),.vcount(vcount), .color(erode), .pixel(eroded));
	////erosion
	//assign black_white = (switch[3])?(switch[2]?b_black_white:g_black_white):switch[1]?r_black_white:o_black_white;
	assign black_white = b_black_white+g_black_white+r_black_white+o_black_white;
	///////////
	////////////
	///dialate dlt(.clk(clk), .vclk(tv_in_line_clock1), .fvh(fvh), .dv(dv), .pixel(black_white), .d_pixel(dialated));
	//erode erdd(.clk(clk),.hcount(hcount),.vcount(vcount), .pixel(vr_pixel[7:0]), .color(eroded));
	///////////
   // for storage, take highest-order RGB bits
	
	 //displaying a blob for 
	 
	 wire [10:0] c_x, cx, q1_x, q2_x, q3_x, q4_x;
	 wire [9:0] c_y, cy, q1_y, q2_y, q3_y, q4_y;
	 wire high_data, high_data1;
	 wire [31:0] sum_x, sum_y, white_count, x, y;
	 //centroid cntrd(clk, tv_in_line_clock1, fvh, dv, black_white, c_x, c_y);
    //////// START centroid calcultations
	 ////////
	 wire [10:0] rc1_x, rc2_x, rc3_x, rc4_x;
	 wire [9:0] rc1_y, rc2_y, rc3_y, rc4_y;
	 ////////
	 
	 ///calculate the center of mass of white color 
	 get_centroid gctr(.clk(clk), .vclk(tv_in_line_clock1), .fvh(fvh), .dv(dv),._x(0), ._y(0), .bound(0),.h(0),.w(0), .pixel(black_white), .cx(c_x), .cy(c_y));
	 
	 get_centroid gctr1(.clk(clk), .vclk(tv_in_line_clock1), .fvh(fvh), .dv(dv),._x(c_x), ._y(c_y), .bound(3'b1),.h(200),.w(200), .pixel(black_white), .cx(cx), .cy(cy));
	 //calculate the centers of the corners 
	 get_centroid gctr2(.clk(clk), .vclk(tv_in_line_clock1), .fvh(fvh), .dv(dv),._x(cx), ._y(cy), .bound(3'b10),.h(0),.w(0), .pixel(b_black_white), .cx(rc1_x), .cy(rc1_y));
	 get_centroid gctr3(.clk(clk), .vclk(tv_in_line_clock1), .fvh(fvh), .dv(dv),._x(cx), ._y(cy), .bound(3'b11),.h(0),.w(0), .pixel(b_black_white), .cx(rc2_x), .cy(rc2_y));
	 get_centroid gctr4(.clk(clk), .vclk(tv_in_line_clock1), .fvh(fvh), .dv(dv),._x(cx), ._y(cy), .bound(3'b100), .h(0),.w(0),.pixel(b_black_white), .cx(rc3_x), .cy(rc3_y));
	 get_centroid gctr5(.clk(clk), .vclk(tv_in_line_clock1), .fvh(fvh), .dv(dv),._x(cx), ._y(cy), .bound(3'b101), .h(0),.w(0),.pixel(b_black_white), .cx(rc4_x), .cy(rc4_y));
	 
	 wire [9:0] h1,h2,h3,h4, w1,w2,w3,w4;
	 assign h1 = (cy>rc1_y)?(cy-rc1_y):(rc1_y-cy);
	 assign h2 = (cy>rc2_y)?(cy-rc2_y):(rc2_y-cy);
	 assign h3 = (cy>rc3_y)?(cy-rc3_y):(rc3_y-cy);
	 assign h4 = (cy>rc4_y)?(cy-rc4_y):(rc4_y-cy);
	 
	 assign w1 = (cx>rc1_x)?(cx-rc1_x):(rc1_x-cx);
	 assign w2 = (cx>rc2_x)?(cx-rc2_x):(rc2_x-cx);
	 assign w3 = (cx>rc3_x)?(cx-rc3_x):(rc3_x-cx);
	 assign w4 = (cx>rc4_x)?(cx-rc4_x):(rc4_x-cx);
	 
	 //HERE we recalculate the centers of the corners
	 get_centroid gctra(.clk(clk), .vclk(tv_in_line_clock1), .fvh(fvh), .dv(dv),._x(rc1_x), ._y(rc1_y), .bound(3'b1),.h(h1),.w(w1), .pixel(b_black_white), .cx(q1_x), .cy(q1_y));
	 get_centroid gctrb(.clk(clk), .vclk(tv_in_line_clock1), .fvh(fvh), .dv(dv),._x(rc2_x), ._y(rc2_y), .bound(3'b1),.h(h2),.w(w2), .pixel(b_black_white), .cx(q2_x), .cy(q2_y));
	 get_centroid gctrc(.clk(clk), .vclk(tv_in_line_clock1), .fvh(fvh), .dv(dv),._x(rc3_x), ._y(rc3_y), .bound(3'b1),.h(h3),.w(w3), .pixel(b_black_white), .cx(q3_x), .cy(q3_y));
	 get_centroid gctrd(.clk(clk), .vclk(tv_in_line_clock1), .fvh(fvh), .dv(dv),._x(rc4_x), ._y(rc4_y), .bound(3'b1),.h(h4),.w(w4), .pixel(b_black_white), .cx(q4_x), .cy(q4_y));
	 ////END of centroid calculations 
	 
	 /////START height and width calculations
	 wire [11:0] height1, height2, width1, width2, width0;
	 wire [12:0] t_height,t_width;
	 dist distw0(.clk(clk), .x_start(23), .x_end(89), .y_start(12), .y_end(90), .distance(width0));
	 dist distw1(.clk(clk), .x_start(q1_x), .x_end(q2_x), .y_start(q1_y), .y_end(q2_y), .distance(width1));
	 dist distw2(.clk(clk), .x_start(q3_x), .x_end(q4_x), .y_start(q3_y), .y_end(q4_y), .distance(width2));
	 dist disth1(.clk(clk), .x_start(q3_x), .x_end(q2_x), .y_start(q3_y), .y_end(q2_y), .distance(height1));
	 dist disth2(.clk(clk), .x_start(q1_x), .x_end(q4_x), .y_start(q1_y), .y_end(q4_y), .distance(height2));
	 wire [12:0] half_width1,half_width2,half_height1,half_height2;
    assign 	half_height1 = (height1>>1);
	 assign 	half_height2 = (height2>>1);
	 assign 	half_width1 = (width1>>1);
	 assign 	half_width2 = (width2>>1);
	 
	 assign t_height = half_height1+half_height2;
	 assign t_width =half_width1+ half_width2;
	 //////END of height and with calculations
	 reg [12:0] tf_x, tf_y;
	 reg [10:0] inf_x;
	 reg [9:0] inf_y;
	 
	 always @(posedge clk)begin//centering the pose
	   inf_x<=(cx<=525)?(525-cx):cx;
		inf_y<=(cy<=525)?(525-cy):cy;
	 end 
	 
	 wire [12:0] cntr_x, cntr_y;
	 transform trfm(.clk(clk), .t_height(t_height), .t_width(t_width), .x(inf_x), .y(inf_y), .cv_x(cntr_x), .cv_y(cntr_y));
	 /////END of coordinate transform  
	 //center_calc cenc(.clk(clk),.inframe(in_frame),.hcount(hcount), .vcount(vcount), .pixel(black_white), .cx(cx),.cy(cy));
	 
	 //////IR transmitter
	 reg [10:0] cent_x;
	 reg [9:0] cent_y;
	 
	 always @(posedge clk) begin 
	    cent_x = (switch[1])?(inf_x):(cntr_x>1023)?1536:cntr_x[10:0];
		 cent_y = (switch[1])?(inf_y):(cntr_y>767)?896:cntr_y[9:0];
	 end 
	 
	 wire [2:0] ir_state;
    ir_transmitter irt (.clock(clock_27mhz), .reset(reset), .trigger(trigger), .clear(clear), .x(cent_x), .y(cent_y), 
         .transmit(clear|trigger), .signal_out(user3[31]), .sstate(ir_state));
	 ///////END of IR Transmitter
	 
	 /////START find shape
	 wire [7:0] q_pixel, q1_pixel, q2_pixel, q3_pixel, q4_pixel;
	 
	 get_shape sh(clk, hcount, q1_x, q2_x, vcount, q1_y, q2_y, q1_pixel);
	 get_shape sh1(clk, hcount, q1_x, q4_x, vcount, q1_y, q4_y, q2_pixel);
	 get_shape sh2(clk, hcount, q3_x, q2_x, vcount, q3_y, q2_y, q3_pixel);
	 get_shape s3(clk, hcount, q3_x, q4_x, vcount, q3_y, q4_y, q4_pixel);
	 
	 assign q_pixel = q1_pixel+q2_pixel+q3_pixel+q4_pixel;
	 /////END find shape
	 
	 /////START blob displays 
	 wire [7:0] c_pixel,c1_pixel,c2_pixel,c3_pixel,c4_pixel,c5_pixel,c6_pixel;
	 centroid_disp  yr1(reset, clk, hcount, vcount, cx, cy, c1_pixel);
	 centroid_disp  yr6(reset, clk, hcount, vcount, q1_x, q1_y, c2_pixel);
	 centroid_disp  yr3(reset, clk, hcount, vcount, q2_x, q2_y, c3_pixel);
	 centroid_disp  yr4(reset, clk, hcount, vcount, q3_x, q3_y, c4_pixel);
	 centroid_disp  yr5(reset, clk, hcount, vcount, q4_x, q4_y, c5_pixel);
	 //centroid_disp #(.HEIGHT(50),.WIDTH(50)) yr7(reset, clk, hcount, vcount, cent_x, cent_y, c6_pixel);
	 assign c_pixel = c1_pixel+c2_pixel+c3_pixel+c4_pixel+c5_pixel;//+c6_pixel;
	 ////////END display modules 
	 
	 
   wire [17:0] RGB_trunc;
	/// Tracking Area 
	wire [9:0] height;
	wire [10:0] width;
	//track tr(.clk(clk), .vclk(tv_in_line_clock1), .reset(reset), .fvh(fvh), .dv(dv), .pixel(black_white), .cx(cx), .cy(cy), .height(height), .width(width));
	wire [7:0] box_pixel;
	assign box_pixel = 0;
	//bounding_box box(.clock(clk), .params(0),.hcount(hcount), .width(width),.x(cx), .vcount(vcount), .height(height),.y(cy), .pixel(box_pixel));
   //assign RGB_trunc = {R[7:2], G[7:2], B[7:2]};
	assign RGB_trunc = (switch[2])?{dialated[7:2], dialated[7:2], dialated[7:2]}:(switch[5])?{R[7:2], G[7:2], B[7:2]}:{black_white[7:2],black_white[7:2],black_white[7:2]};

   // code to write NTSC data to video memory

   wire [18:0] ntsc_addr;
   wire [35:0] ntsc_data;
   wire        ntsc_we;
   ntsc_to_zbt n2z (clk, tv_in_line_clock1, fvh, dv, RGB_trunc,
		    ntsc_addr, ntsc_data, ntsc_we, switch[6]);//{_rgb[23:18], _rgb[15:9], _rgb[7:2]}

   // code to write pattern to ZBT memory
   reg [31:0] 	count;
   always @(posedge clk) count <= reset ? 0 : count + 1;

   wire [18:0] 	vram_addr2 = count[0+18:0];
   wire [35:0] 	vpat = ( switch[1] ? {4{count[3+3:3],4'b0}}
			 : {4{count[3+4:4],4'b0}} );

   // mux selecting read/write to memory based on which write-enable is chosen

   wire 	sw_ntsc = ~switch[7];
//   wire 	my_we = sw_ntsc ? (hcount[1:0]==2'd2) : blank;
   wire 	my_we = sw_ntsc ? hcount[0] : blank;
   wire [18:0] 	write_addr = sw_ntsc ? ntsc_addr : vram_addr2;
   wire [35:0] 	write_data = sw_ntsc ? ntsc_data : vpat;

//   wire 	write_enable = sw_ntsc ? (my_we & ntsc_we) : my_we;
//   assign 	vram_addr = write_enable ? write_addr : vram_addr1;
//   assign 	vram_we = write_enable;

   assign 	vram_addr = my_we ? write_addr : vram_addr1;
   assign 	vram_we = my_we;
   assign 	vram_write_data = write_data;

   // select output pixel data

   reg [17:0] 	pixel;
   reg 	b,hs,vs;
   
	//wire [10:0] out;
   //sqrt_func sqrt(cx, out, clk);	

   always @(posedge clk)
     begin
	pixel <= (q_pixel==8'hFF)?{12'b0, q_pixel[7:2]}:((box_pixel==8'hFF)?{box_pixel[7:2], 12'b0}:(switch[4])?(vr_pixel[7:2]<=c_pixel[7:2])?{c_pixel[7:2], c_pixel[7:2], c_pixel[7:2]}:vr_pixel:(switch[0] ? {hcount[8:6],15'b0} : vr_pixel));
	b <= blank;
	hs <= hsync;
	vs <= vsync;
     end
/*
   assign pixel = vr_pixel;
   delayN #(.NDELAY(3)) b_delay(clk, blank, b);
   delayN #(.NDELAY(3)) h_delay(clk, hsync, hs);
   delayN #(.NDELAY(3)) v_delay(clk, vsync, vs);
*/

   // Video filter module for each pixel
   

   // VGA Output.  In order to meet the setup and hold times of the
   // AD7125, we send it ~clk.
    //wire [21:0] sum_sq;
	 //assign sum_sq = 4100;
	 //wire [10:0]  x_out;
    //sqrt_func sqrt1(.x_in(sum_sq), .clk(clk), .x_out(x_out), .rdy(rdy) );
   //assign vga_out_red = pixel_filtered[23:16];
   //assign vga_out_green = pixel_filtered[15:8];
   //assign vga_out_blue = pixel_filtered[7:0];

   assign vga_out_red =  {pixel[17:12], 2'b0};
   assign vga_out_green = {pixel[11:6], 2'b0};
   assign vga_out_blue = {pixel[5:0], 2'b0};

   assign vga_out_sync_b = 1'b1;    // not used
   assign vga_out_pixel_clock = ~clk;
   assign vga_out_blank_b = ~b;
   assign vga_out_hsync = hs;
   assign vga_out_vsync = vs;

   // debugging
   wire [12:0] disp_x, disp_y;
	assign disp_x = (switch[0])?{2'b0, cx}:cntr_x;
	assign disp_y = (switch[0])?{3'b0, cy}:cntr_y;
	
   assign led = ~{vram_addr[18:12],white,reseted,divided};
   assign analyzer3_data = {8'b0, 4'b0,tv_in_line_clock1,fvh};
	assign analyzer3_clock = tv_in_line_clock1;
   always @(posedge clk)
     // dispdata <= {vram_read_data,9'b0,vram_addr};
     //dispdata <= {ntsc_data,1'b0,fvh,3'b0,c_x,c_y,2'b0};
	  
	  dispdata <= {disp_x,4'b0, disp_y, t_width, t_height,5'b0,ir_state};

	
endmodule


///////////////////////////////////////////////////////////////////////////////
// xvga: Generate XVGA display signals (1024 x 768 @ 60Hz)

module xvga(vclock,hcount,vcount,hsync,vsync,blank);
   input vclock;
   output [10:0] hcount;
   output [9:0] vcount;
   output 	vsync;
   output 	hsync;
   output 	blank;

   reg 	  hsync,vsync,hblank,vblank,blank;
   reg [10:0] 	 hcount;    // pixel number on current line
   reg [9:0] vcount;	 // line number

   // horizontal: 1344 pixels total
   // display 1024 pixels per line
   wire      hsyncon,hsyncoff,hreset,hblankon;
   assign    hblankon = (hcount == 1023);    
   assign    hsyncon = (hcount == 1047);
   assign    hsyncoff = (hcount == 1183);
   assign    hreset = (hcount == 1343);

   // vertical: 806 lines total
   // display 768 lines
   wire      vsyncon,vsyncoff,vreset,vblankon;
   assign    vblankon = hreset & (vcount == 767);    
   assign    vsyncon = hreset & (vcount == 776);
   assign    vsyncoff = hreset & (vcount == 782);
   assign    vreset = hreset & (vcount == 805);

   // sync and blanking
   wire      next_hblank,next_vblank;
   assign next_hblank = hreset ? 0 : hblankon ? 1 : hblank;
   assign next_vblank = vreset ? 0 : vblankon ? 1 : vblank;
   always @(posedge vclock) begin
      hcount <= hreset ? 0 : hcount + 1;
      hblank <= next_hblank;
      hsync <= hsyncon ? 0 : hsyncoff ? 1 : hsync;  // active low

      vcount <= hreset ? (vreset ? 0 : vcount + 1) : vcount;
      vblank <= next_vblank;
      vsync <= vsyncon ? 0 : vsyncoff ? 1 : vsync;  // active low

      blank <= next_vblank | (next_hblank & ~hreset);
   end
endmodule


module vram_display(reset,clk,hcount,vcount,vr_pixel,center_x, center_y, hold_count, hold_x, hold_y, reseted, divided,white,
		    vram_addr,vram_read_data);

   input reset, clk;
   input [10:0] hcount;
   input [9:0] 	vcount;
   output [17:0] vr_pixel;
   output [18:0] vram_addr;
   input [35:0]  vram_read_data;
	
	output reg [10:0] center_x;
	output reg [9:0] center_y;
	
	output reg divided, reseted;
	output white;
	output reg [31:0]  hold_x, hold_y, hold_count;
	////accumulation registers 
	reg [32:0] sum_x;
	reg [32:0] sum_y;
	reg [31:0] white_count;

   //forecast hcount & vcount 8 clock cycles ahead to get data from ZBT
   wire [10:0] hcount_f = (hcount >= 1048) ? (hcount - 1048) : (hcount + 8);
   wire [9:0] vcount_f = (hcount >= 1048) ? ((vcount == 805) ? 0 : vcount + 1) : vcount;
      
   wire [18:0] 	 vram_addr = {vcount_f, hcount_f[9:1]};


//   wire [1:0] 	 hc4 = hcount[1:0];
   wire [1:0] hc2 = hcount[0];
   reg [17:0] 	 vr_pixel;
   reg [35:0] 	 vr_data_latched;
   reg [35:0] 	 last_vr_data;
	
   //division registers
	
	wire [31:0] quot_x, quot_y,rem_x, rem_y; 
	wire x_rdy, y_rdy;
	

/*
   always @(posedge clk)
     last_vr_data <= (hc4==2'd3) ? vr_data_latched : last_vr_data;
   always @(posedge clk)
     vr_data_latched <= (hc4==2'd1) ? vram_read_data : vr_data_latched;
   always @(*)		// each 36-bit word from RAM is decoded to 4 bytes
     case (hc4)
       2'd3: vr_pixel = last_vr_data[7:0];
       2'd2: vr_pixel = last_vr_data[7+8:0+8];
       2'd1: vr_pixel = last_vr_data[7+16:0+16];
       2'd0: vr_pixel = last_vr_data[7+24:0+24];
     endcase
*/
   wire rst = (hcount==0 & vcount==0);
	wire divide = ((hcount==0) & (vcount==767));//
	
	//assign reseted=(rst)?~reseted:reseted;
	//assign divided = (divide)?~divided:divided;
	always @(*) begin 
		reseted=(rst)?~reseted:reseted;
	   divided = (divide)?~divided:divided;
	end
// Modification for color
   always @(posedge clk)
     last_vr_data <= (hc2) ? vr_data_latched : last_vr_data;

   always @(posedge clk)
     vr_data_latched <= (~hc2) ? vram_read_data : vr_data_latched;
   assign white  = (last_vr_data[17:10]>30);
   always @(*)		// each 36-bit word from RAM is decoded to 4 bytes
     case (hc2)
       1'd1: begin vr_pixel = last_vr_data[17:0];
				sum_x=(rst)?0:(last_vr_data[17:10]>30)?sum_x+hcount: sum_x;
				sum_y=(rst)?0:(last_vr_data[17:10]>30)?sum_y+vcount: sum_y;
				white_count=(rst)?0:(last_vr_data[17:10]>30)?white_count+1: white_count;
			end 
       1'd0: begin vr_pixel = last_vr_data[35:18];
				sum_x=(rst)?0:(last_vr_data[35:30]>30)?sum_x+hcount: sum_x;
				sum_y=(rst)?0:(last_vr_data[35:30]>30)?sum_y+vcount: sum_y;
				white_count=(rst)?0:(last_vr_data[35:30]>30)?white_count+1: white_count;
				end
     endcase
	always @(posedge clk) begin 
	     hold_x=(divide)?sum_x: hold_x;
		  hold_y=(divide)?sum_y: hold_y;
		  hold_count=(divide)?white_count: hold_count;
		  
		  center_x = (x_rdy)?quot_x[10:0]: center_x;
		  center_y = (x_rdy)?quot_y[9:0]: center_y;
	end 
	_divider #(.WIDTH(32)) 
  div1(.clk(clk), .sign(0), .start(divide),.dividend(hold_x), .divisor(hold_count),.quotient(quot_x),.remainder(rem_x),.ready(x_rdy));
  _divider #(.WIDTH(32)) 
  div2(.clk(clk), .sign(0), .start(divide),.dividend(hold_y), .divisor(hold_count),.quotient(quot_y),.remainder(rem_y),.ready(y_rdy));

endmodule // vram_display

/////////////////////////////////////////////////////////////////////////////
// parameterized delay line 

module delayN(clk,in,out);
   input clk;
   input in;
   output out;

   parameter NDELAY = 3;

   reg [NDELAY-1:0] shiftreg;
   wire 	    out = shiftreg[NDELAY-1];

   always @(posedge clk)
     shiftreg <= {shiftreg[NDELAY-2:0],in};

endmodule // delayN

////////////////////////////////////////////////////////////////////////////
// ramclock module

///////////////////////////////////////////////////////////////////////////////
//
// 6.111 FPGA Labkit -- ZBT RAM clock generation
//
//
// Created: April 27, 2004
// Author: Nathan Ickes
//
///////////////////////////////////////////////////////////////////////////////
//
// This module generates deskewed clocks for driving the ZBT SRAMs and FPGA 
// registers. A special feedback trace on the labkit PCB (which is length 
// matched to the RAM traces) is used to adjust the RAM clock phase so that 
// rising clock edges reach the RAMs at exactly the same time as rising clock 
// edges reach the registers in the FPGA.
//
// The RAM clock signals are driven by DDR output buffers, which further 
// ensures that the clock-to-pad delay is the same for the RAM clocks as it is 
// for any other registered RAM signal.
//
// When the FPGA is configured, the DCMs are enabled before the chip-level I/O
// drivers are released from tristate. It is therefore necessary to
// artificially hold the DCMs in reset for a few cycles after configuration. 
// This is done using a 16-bit shift register. When the DCMs have locked, the 
// <lock> output of this mnodule will go high. Until the DCMs are locked, the 
// ouput clock timings are not guaranteed, so any logic driven by the 
// <fpga_clock> should probably be held inreset until <locked> is high.
//
///////////////////////////////////////////////////////////////////////////////

module ramclock(ref_clock, fpga_clock, ram0_clock, ram1_clock, 
	        clock_feedback_in, clock_feedback_out, locked);
   
   input ref_clock;                 // Reference clock input
   output fpga_clock;               // Output clock to drive FPGA logic
   output ram0_clock, ram1_clock;   // Output clocks for each RAM chip
   input  clock_feedback_in;        // Output to feedback trace
   output clock_feedback_out;       // Input from feedback trace
   output locked;                   // Indicates that clock outputs are stable
   
   wire  ref_clk, fpga_clk, ram_clk, fb_clk, lock1, lock2, dcm_reset;

   ////////////////////////////////////////////////////////////////////////////
   
   //To force ISE to compile the ramclock, this line has to be removed.
   //IBUFG ref_buf (.O(ref_clk), .I(ref_clock));
	
	assign ref_clk = ref_clock;
   
   BUFG int_buf (.O(fpga_clock), .I(fpga_clk));

   DCM int_dcm (.CLKFB(fpga_clock),
		.CLKIN(ref_clk),
		.RST(dcm_reset),
		.CLK0(fpga_clk),
		.LOCKED(lock1));
   // synthesis attribute DLL_FREQUENCY_MODE of int_dcm is "LOW"
   // synthesis attribute DUTY_CYCLE_CORRECTION of int_dcm is "TRUE"
   // synthesis attribute STARTUP_WAIT of int_dcm is "FALSE"
   // synthesis attribute DFS_FREQUENCY_MODE of int_dcm is "LOW"
   // synthesis attribute CLK_FEEDBACK of int_dcm  is "1X"
   // synthesis attribute CLKOUT_PHASE_SHIFT of int_dcm is "NONE"
   // synthesis attribute PHASE_SHIFT of int_dcm is 0
   
   BUFG ext_buf (.O(ram_clock), .I(ram_clk));
   
   IBUFG fb_buf (.O(fb_clk), .I(clock_feedback_in));
   
   DCM ext_dcm (.CLKFB(fb_clk), 
		    .CLKIN(ref_clk), 
		    .RST(dcm_reset),
		    .CLK0(ram_clk),
		    .LOCKED(lock2));
   // synthesis attribute DLL_FREQUENCY_MODE of ext_dcm is "LOW"
   // synthesis attribute DUTY_CYCLE_CORRECTION of ext_dcm is "TRUE"
   // synthesis attribute STARTUP_WAIT of ext_dcm is "FALSE"
   // synthesis attribute DFS_FREQUENCY_MODE of ext_dcm is "LOW"
   // synthesis attribute CLK_FEEDBACK of ext_dcm  is "1X"
   // synthesis attribute CLKOUT_PHASE_SHIFT of ext_dcm is "NONE"
   // synthesis attribute PHASE_SHIFT of ext_dcm is 0

   SRL16 dcm_rst_sr (.D(1'b0), .CLK(ref_clk), .Q(dcm_reset),
		     .A0(1'b1), .A1(1'b1), .A2(1'b1), .A3(1'b1));
   // synthesis attribute init of dcm_rst_sr is "000F";
   

   OFDDRRSE ddr_reg0 (.Q(ram0_clock), .C0(ram_clock), .C1(~ram_clock),
		      .CE (1'b1), .D0(1'b1), .D1(1'b0), .R(1'b0), .S(1'b0));
   OFDDRRSE ddr_reg1 (.Q(ram1_clock), .C0(ram_clock), .C1(~ram_clock),
		      .CE (1'b1), .D0(1'b1), .D1(1'b0), .R(1'b0), .S(1'b0));
   OFDDRRSE ddr_reg2 (.Q(clock_feedback_out), .C0(ram_clock), .C1(~ram_clock),
		      .CE (1'b1), .D0(1'b1), .D1(1'b0), .R(1'b0), .S(1'b0));

   assign locked = lock1 && lock2;
   
endmodule


