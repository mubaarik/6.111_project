///////////////////////////////////////////////////////////////////////////////
//
// Pushbutton Debounce Module (video version - 24 bits)  
//
///////////////////////////////////////////////////////////////////////////////

module debounce (input reset, clock, noisy,output reg clean);

   reg [19:0] count;
   reg new;

   always @(posedge clock)
     if (reset) begin new <= noisy; clean <= noisy; count <= 0; end
     else if (noisy != new) begin new <= noisy; count <= 0; end
     else if (count == 650000) clean <= new;
     else count <= count+1;

endmodule

///////////////////////////////////////////////////////////////////////////////
//
// 6.111 FPGA Labkit -- Template Toplevel Module
//
// For Labkit Revision 004
//
//
// Created: October 31, 2004, from revision 003 file
// Author: Nathan Ickes
//
///////////////////////////////////////////////////////////////////////////////
//
// CHANGES FOR BOARD REVISION 004
//
// 1) Added signals for logic analyzer pods 2-4.
// 2) Expanded "tv_in_ycrcb" to 20 bits.
// 3) Renamed "tv_out_data" to "tv_out_i2c_data" and "tv_out_sclk" to
//    "tv_out_i2c_clock".
// 4) Reversed disp_data_in and disp_data_out signals, so that "out" is an
//    output of the FPGA, and "in" is an input.
//
// CHANGES FOR BOARD REVISION 003
//
// 1) Combined flash chip enables into a single signal, flash_ce_b.
//
// CHANGES FOR BOARD REVISION 002
//
// 1) Added SRAM clock feedback path input and output
// 2) Renamed "mousedata" to "mouse_data"
// 3) Renamed some ZBT memory signals. Parity bits are now incorporated into 
//    the data bus, and the byte write enables have been combined into the
//    4-bit ram#_bwe_b bus.
// 4) Removed the "systemace_clock" net, since the SystemACE clock is now
//    hardwired on the PCB to the oscillator.
//
///////////////////////////////////////////////////////////////////////////////
//
// Complete change history (including bug fixes)
//
// 2012-Sep-15: Converted to 24bit RGB
//
// 2005-Sep-09: Added missing default assignments to "ac97_sdata_out",
//              "disp_data_out", "analyzer[2-3]_clock" and
//              "analyzer[2-3]_data".
//
// 2005-Jan-23: Reduced flash address bus to 24 bits, to match 128Mb devices
//              actually populated on the boards. (The boards support up to
//              256Mb devices, with 25 address lines.)
//
// 2004-Oct-31: Adapted to new revision 004 board.
//
// 2004-May-01: Changed "disp_data_in" to be an output, and gave it a default
//              value. (Previous versions of this file declared this port to
//              be an input.)
///
// 2004-Apr-29: Reduced SRAM address busses to 19 bits, to match 18Mb devices
//              actually populated on the boards. (The boards support up to
//              72Mb devices, with 21 address lines.)
//
// 2004-Apr-29: Change history started
//
///////////////////////////////////////////////////////////////////////////////

module lab3   (beep, audio_reset_b, ac97_sdata_out, ac97_sdata_in, ac97_synch,
	       ac97_bit_clock,
	       
	       vga_out_red, vga_out_green, vga_out_blue, vga_out_sync_b,
	       vga_out_blank_b, vga_out_pixel_clock, vga_out_hsync,
	       vga_out_vsync,

	       tv_out_ycrcb, tv_out_reset_b, tv_out_clock, tv_out_i2c_clock,
	       tv_out_i2c_data, tv_out_pal_ntsc, tv_out_hsync_b,
	       tv_out_vsync_b, tv_out_blank_b, tv_out_subcar_reset,

	       tv_in_ycrcb, tv_in_data_valid, tv_in_line_clock1,
	       tv_in_line_clock2, tv_in_aef, tv_in_hff, tv_in_aff,
	       tv_in_i2c_clock, tv_in_i2c_data, tv_in_fifo_read,
	       tv_in_fifo_clock, tv_in_iso, tv_in_reset_b, tv_in_clock,

	       ram0_data, ram0_address, ram0_adv_ld, ram0_clk, ram0_cen_b,
	       ram0_ce_b, ram0_oe_b, ram0_we_b, ram0_bwe_b, 

	       ram1_data, ram1_address, ram1_adv_ld, ram1_clk, ram1_cen_b,
	       ram1_ce_b, ram1_oe_b, ram1_we_b, ram1_bwe_b,

	       clock_feedback_out, clock_feedback_in,

	       flash_data, flash_address, flash_ce_b, flash_oe_b, flash_we_b,
	       flash_reset_b, flash_sts, flash_byte_b,

	       rs232_txd, rs232_rxd, rs232_rts, rs232_cts,

	       mouse_clock, mouse_data, keyboard_clock, keyboard_data,

	       clock_27mhz, clock1, clock2,

	       disp_blank, disp_data_out, disp_clock, disp_rs, disp_ce_b,
	       disp_reset_b, disp_data_in,

	       button0, button1, button2, button3, button_enter, button_right,
	       button_left, button_down, button_up,

	       switch,

	       led,
	       
	       user1, user2, user3, user4,
	       
	       daughtercard,

	       systemace_data, systemace_address, systemace_ce_b,
	       systemace_we_b, systemace_oe_b, systemace_irq, systemace_mpbrdy,
	       
	       analyzer1_data, analyzer1_clock,
 	       analyzer2_data, analyzer2_clock,
 	       analyzer3_data, analyzer3_clock,
 	       analyzer4_data, analyzer4_clock);

   output beep, audio_reset_b, ac97_synch, ac97_sdata_out;
   input  ac97_bit_clock, ac97_sdata_in;
   
   output [7:0] vga_out_red, vga_out_green, vga_out_blue;
   output vga_out_sync_b, vga_out_blank_b, vga_out_pixel_clock,
	  vga_out_hsync, vga_out_vsync;

   output [9:0] tv_out_ycrcb;
   output tv_out_reset_b, tv_out_clock, tv_out_i2c_clock, tv_out_i2c_data,
	  tv_out_pal_ntsc, tv_out_hsync_b, tv_out_vsync_b, tv_out_blank_b,
	  tv_out_subcar_reset;
   
   input  [19:0] tv_in_ycrcb;
   input  tv_in_data_valid, tv_in_line_clock1, tv_in_line_clock2, tv_in_aef,
	  tv_in_hff, tv_in_aff;
   output tv_in_i2c_clock, tv_in_fifo_read, tv_in_fifo_clock, tv_in_iso,
	  tv_in_reset_b, tv_in_clock;
   inout  tv_in_i2c_data;
        
   inout  [35:0] ram0_data;
   output [18:0] ram0_address;
   output ram0_adv_ld, ram0_clk, ram0_cen_b, ram0_ce_b, ram0_oe_b, ram0_we_b;
   output [3:0] ram0_bwe_b;
   
   inout  [35:0] ram1_data;
   output [18:0] ram1_address;
   output ram1_adv_ld, ram1_clk, ram1_cen_b, ram1_ce_b, ram1_oe_b, ram1_we_b;
   output [3:0] ram1_bwe_b;

   input  clock_feedback_in;
   output clock_feedback_out;
   
   inout  [15:0] flash_data;
   output [24:0] flash_address;
   output flash_ce_b, flash_oe_b, flash_we_b, flash_reset_b, flash_byte_b;
   input  flash_sts;
   
   output rs232_txd, rs232_rts;
   input  rs232_rxd, rs232_cts;

   input  mouse_clock, mouse_data, keyboard_clock, keyboard_data;

   input  clock_27mhz, clock1, clock2;

   output disp_blank, disp_clock, disp_rs, disp_ce_b, disp_reset_b;  
   input  disp_data_in;
   output  disp_data_out;
   
   input  button0, button1, button2, button3, button_enter, button_right,
	  button_left, button_down, button_up;
   input  [7:0] switch;
   output [7:0] led;

   inout [31:0] user1, user2, user3, user4;
   
   inout [43:0] daughtercard;

   inout  [15:0] systemace_data;
   output [6:0]  systemace_address;
   output systemace_ce_b, systemace_we_b, systemace_oe_b;
   input  systemace_irq, systemace_mpbrdy;

   output [15:0] analyzer1_data, analyzer2_data, analyzer3_data, 
		 analyzer4_data;
   output analyzer1_clock, analyzer2_clock, analyzer3_clock, analyzer4_clock;

   ////////////////////////////////////////////////////////////////////////////
   //
   // I/O Assignments
   //
   ////////////////////////////////////////////////////////////////////////////
   
   // Audio Input and Output
   assign beep= 1'b0;
   //assign audio_reset_b = 1'b0;
   //assign ac97_synch = 1'b0;
   //assign ac97_sdata_out = 1'b0;
   // ac97_sdata_in is an input

   // Video Output
   assign tv_out_ycrcb = 10'h0;
   assign tv_out_reset_b = 1'b0;
   assign tv_out_clock = 1'b0;
   assign tv_out_i2c_clock = 1'b0;
   assign tv_out_i2c_data = 1'b0;
   assign tv_out_pal_ntsc = 1'b0;
   assign tv_out_hsync_b = 1'b1;
   assign tv_out_vsync_b = 1'b1;
   assign tv_out_blank_b = 1'b1;
   assign tv_out_subcar_reset = 1'b0;
   
   // Video Input
   assign tv_in_i2c_clock = 1'b0;
   assign tv_in_fifo_read = 1'b0;
   assign tv_in_fifo_clock = 1'b0;
   assign tv_in_iso = 1'b0;
   assign tv_in_reset_b = 1'b0;
   assign tv_in_clock = 1'b0;
   assign tv_in_i2c_data = 1'bZ;
   // tv_in_ycrcb, tv_in_data_valid, tv_in_line_clock1, tv_in_line_clock2, 
   // tv_in_aef, tv_in_hff, and tv_in_aff are inputs
   
   // SRAMs
   assign ram0_data = 36'hZ;
   assign ram0_address = 19'h0;
   assign ram0_adv_ld = 1'b0;
   assign ram0_clk = 1'b0;
   assign ram0_cen_b = 1'b1;
   assign ram0_ce_b = 1'b1;
   assign ram0_oe_b = 1'b1;
   assign ram0_we_b = 1'b1;
   assign ram0_bwe_b = 4'hF;
   assign ram1_data = 36'hZ; 
   assign ram1_address = 19'h0;
   assign ram1_adv_ld = 1'b0;
   assign ram1_clk = 1'b0;
   assign ram1_cen_b = 1'b1;
   assign ram1_ce_b = 1'b1;
   assign ram1_oe_b = 1'b1;
   assign ram1_we_b = 1'b1;
   assign ram1_bwe_b = 4'hF;
   assign clock_feedback_out = 1'b0;
   // clock_feedback_in is an input
   
   // Flash ROM
   assign flash_data = 16'hZ;
   assign flash_address = 25'h0;
   assign flash_ce_b = 1'b1;
   assign flash_oe_b = 1'b1;
   assign flash_we_b = 1'b1;
   assign flash_reset_b = 1'b0;
   assign flash_byte_b = 1'b1;
   // flash_sts is an input

   // RS-232 Interface
   assign rs232_txd = 1'b1;
   assign rs232_rts = 1'b1;
   // rs232_rxd and rs232_cts are inputs

   // PS/2 Ports
   // mouse_clock, mouse_data, keyboard_clock, and keyboard_data are inputs

   // LED Displays
   //assign disp_blank = 1'b1;
//   assign disp_clock = 1'b0;
//   assign disp_rs = 1'b0;
//   assign disp_ce_b = 1'b1;
//   assign disp_reset_b = 1'b0;
//   assign disp_data_out = 1'b0;
   // disp_data_in is an input

   // Buttons, Switches, and Individual LEDs
   //lab3 assign led = 8'hFF;
   // button0, button1, button2, button3, button_enter, button_right,
   // button_left, button_down, button_up, and switches are inputs

   // User I/Os
   assign user1 = 32'hZ;
   assign user2 = 32'hZ;
   assign user3 = 32'hZ;
   assign user4 = 32'hZ;

   // Daughtercard Connectors
   assign daughtercard = 44'hZ;

   // SystemACE Microprocessor Port
   assign systemace_data = 16'hZ;
   assign systemace_address = 7'h0;
   assign systemace_ce_b = 1'b1;
   assign systemace_we_b = 1'b1;
   assign systemace_oe_b = 1'b1;
   // systemace_irq and systemace_mpbrdy are inputs

   // Logic Analyzer
   assign analyzer1_data = 16'h0;
   assign analyzer1_clock = 1'b1;
   assign analyzer2_data = 16'h0;
   assign analyzer2_clock = 1'b1;
   assign analyzer3_data = 16'h0;
   assign analyzer3_clock = 1'b1;
   assign analyzer4_data = 16'h0;
   assign analyzer4_clock = 1'b1;
			    
   ////////////////////////////////////////////////////////////////////////////
   //
   // lab3 : a simple pong game
   //
   ////////////////////////////////////////////////////////////////////////////

   // use FPGA's digital clock manager to produce a
   // 65MHz clock (actually 64.8MHz)
   wire clock_65mhz_unbuf,clock_65mhz;
   DCM vclk1(.CLKIN(clock_27mhz),.CLKFX(clock_65mhz_unbuf));
   // synthesis attribute CLKFX_DIVIDE of vclk1 is 10
   // synthesis attribute CLKFX_MULTIPLY of vclk1 is 24
   // synthesis attribute CLK_FEEDBACK of vclk1 is NONE
   // synthesis attribute CLKIN_PERIOD of vclk1 is 37
   BUFG vclk2(.O(clock_65mhz),.I(clock_65mhz_unbuf));

   // power-on reset generation
   wire power_on_reset;    // remain high for first 16 clocks
   SRL16 reset_sr (.D(1'b0), .CLK(clock_65mhz), .Q(power_on_reset),
		   .A0(1'b1), .A1(1'b1), .A2(1'b1), .A3(1'b1));
   defparam reset_sr.INIT = 16'hFFFF;

   // ENTER button is user reset
   wire reset,user_reset;
   debounce db1(.reset(power_on_reset),.clock(clock_65mhz),.noisy(~button0),.clean(user_reset));
   assign reset = user_reset | power_on_reset;


   ///////HERE WE HAVE THE SOUND

             
   wire [7:0] from_ac97_data, to_ac97_data;
   wire ready;

   // allow user to adjust volume
   wire vup,vdown;
   reg old_vup,old_vdown;
   debounce bup(.reset(reset),.clock(clock_27mhz),.noisy(~button_up),.clean(vup));
   debounce bdown(.reset(reset),.clock(clock_27mhz),.noisy(~button_down),.clean(vdown));
   reg [4:0] volume;
   always @ (posedge clock_27mhz) begin
     if (reset) volume <= 5'd8;
     else begin
   if (vup & ~old_vup & volume != 5'd31) volume <= volume+1;       
   if (vdown & ~old_vdown & volume != 5'd0) volume <= volume-1;       
     end
     old_vup <= vup;
     old_vdown <= vdown;
   end

   // AC97 driver
   lab5audio a(clock_27mhz, reset, volume, from_ac97_data, to_ac97_data, ready,
          audio_reset_b, ac97_sdata_out, ac97_sdata_in,
          ac97_synch, ac97_bit_clock);

   // push ENTER button to record, release to playback
   wire trigger, counting;
   wire playback,_trigger;
   //assign _trigger = trigger;
   debounce benter(.reset(reset),.clock(clock_27mhz),.noisy(button_enter),.clean(playback));
   //debounce bu3(.reset(reset),.clock(clock_27mhz),.noisy(~button3),.clean(_trigger));
   // switch 0 up for filtering, down for no filtering
   wire filter;
   debounce sw0(.reset(reset),.clock(clock_27mhz),.noisy(switch[7]),.clean(filter));
   wire echo, move;
   debounce sw1(.reset(reset),.clock(clock_27mhz),.noisy(switch[6]),.clean(echo));
   debounce sw5(.reset(reset),.clock(clock_27mhz),.noisy(switch[5]),.clean(move));
   // light up LEDs when recording, show volume during playback.
   // led is active low
   ///assign led = playback ? ~{filter,button_enter,1'b0, volume} : ~{filter,1'b0,6'hFF};

   // record module
   recorder r(.clock(clock_27mhz), .reset(reset), .ready(ready),
              .playback(playback),.echo(echo),.trigger(_trigger), .filter(filter),
              .from_ac97_data(from_ac97_data),.to_ac97_data(to_ac97_data));
  ////////END OF SOUND STUFF

   
   ////display
	wire [63:0] data;
	display_16hex disppp(reset, clock_27mhz, data, 
		disp_blank, disp_clock, disp_rs, disp_ce_b,
		disp_reset_b, disp_data_out);
   // generate basic XVGA video signals
   wire [10:0] hcount;
   wire [9:0]  vcount;
   wire hsync,vsync,blank;
   xvga xvga1(.vclock(clock_65mhz),.hcount(hcount),.vcount(vcount),
              .hsync(hsync),.vsync(vsync),.blank(blank));

   // feed XVGA signals to user's pong game
	wire sync_serial;
   synchronize s_serial(.clk(clock_27mhz), .in(user3[30]), .out(sync_serial));
	
   wire [23:0] pixel;
   wire phsync,pvsync,pblank;
   wire [10:0] x;
   wire [9:0] y;

   display pg(.vclock(clock_65mhz), .clk(clock_27mhz),.reset(reset), .sync_serial(sync_serial),.move(move),
		.hcount(hcount),.vcount(vcount), .keyboard_clock(keyboard_clock),
                .hsync(hsync),.vsync(vsync),.blank(blank), .keyboard_data(keyboard_data),.have_trigger(_trigger),
		.phsync(phsync),.pvsync(pvsync),.pblank(pblank),.pixel(pixel), ._x(x), ._y(y), 
		.show_trigger(trigger), .counting(counting));
   
	 
	 wire [7:0] c_pixel;
	 
	 //////////
	 
	 //centroid_disp yr1(.reset(reset), .clk(vclock), .hcount(hcount), .vcount(vcount), .x(64), .y(64), .pixel(c_pixel));
   // switch[1:0] selects which video generator to use:
   //  00: user's pong game
   //  01: 1 pixel outline of active video area (adjust screen controls)
   //  10: color bars
   reg [23:0] rgb;
   wire border = (hcount==0 | hcount==1023 | vcount==0 | vcount==767);
   
   reg b,hs,vs;
   always @(posedge clock_65mhz) begin
      if (switch[1:0] == 2'b01) begin
	 // 1 pixel outline of visible area (white)
	 hs <= hsync;
	 vs <= vsync;
	 b <= blank;
	 rgb <= {24{border}};
      end else if (switch[1:0] == 2'b10) begin
	 // color bars
	 hs <= hsync;
	 vs <= vsync;
	 b <= blank;
	 rgb <= {{8{hcount[8]}}, {8{hcount[7]}}, {8{hcount[6]}}} ;
      end else begin
         // default: pong
	 hs <= phsync;
	 vs <= pvsync;
	 b <= pblank;
	 rgb <= (switch[4])?{c_pixel,c_pixel,c_pixel}:pixel;
      end
   end


//////random testing area
wire [11:0] dist;
wire [21:0] sum_sqrs;
dist dist1(.clk(clock_65mhz), .x_start(98), .x_end(198), .y_start(90), .y_end(239), .distance(dist), .sum_sqrs(sum_sqrs));
/////////////
   // VGA Output.  In order to meet the setup and hold times of the
   // AD7125, we send it ~clock_65mhz.
   assign vga_out_red = rgb[23:16];
   assign vga_out_green = rgb[15:8];
   assign vga_out_blue = rgb[7:0];
   assign vga_out_sync_b = 1'b1;    // not used
   assign vga_out_blank_b = ~b;
   assign vga_out_pixel_clock = ~clock_65mhz;
   assign vga_out_hsync = hs;
   assign vga_out_vsync = vs;
   
   assign led = ~{1'b0,~counting,~trigger,reset,switch[1:0]};
   assign data =  {dist, 4'b0, x, 4'b0, y};
endmodule

////////////////////////////////////////////////////////////////////////////////
//
// xvga: Generate XVGA display signals (1024 x 768 @ 60Hz)
//
////////////////////////////////////////////////////////////////////////////////

module xvga(input vclock,
            output reg [10:0] hcount,    // pixel number on current line
            output reg [9:0] vcount,	 // line number
            output reg vsync,hsync,blank);

   // horizontal: 1344 pixels total
   // display 1024 pixels per line
   reg hblank,vblank;
   wire hsyncon,hsyncoff,hreset,hblankon;
   assign hblankon = (hcount == 1023);    
   assign hsyncon = (hcount == 1047);
   assign hsyncoff = (hcount == 1183);
   assign hreset = (hcount == 1343);

   // vertical: 806 lines total
   // display 768 lines
   wire vsyncon,vsyncoff,vreset,vblankon;
   assign vblankon = hreset & (vcount == 767);    
   assign vsyncon = hreset & (vcount == 776);
   assign vsyncoff = hreset & (vcount == 782);
   assign vreset = hreset & (vcount == 805);

   // sync and blanking
   wire next_hblank,next_vblank;
   assign next_hblank = hreset ? 0 : hblankon ? 1 : hblank;
   assign next_vblank = vreset ? 0 : vblankon ? 1 : vblank;
   always @(posedge vclock) begin
      hcount <= hreset ? 0 : hcount + 1;
      hblank <= next_hblank;
      hsync <= hsyncon ? 0 : hsyncoff ? 1 : hsync;  // active low

      vcount <= hreset ? (vreset ? 0 : vcount + 1) : vcount;
      vblank <= next_vblank;
      vsync <= vsyncon ? 0 : vsyncoff ? 1 : vsync;  // active low

      blank <= next_vblank | (next_hblank & ~hreset);
   end
endmodule

////////////////////////////////////////////////////////////////////////////////
//
// pong_game: the game itself!
//
////////////////////////////////////////////////////////////////////////////////

module display (
   input vclock, clk,	// 65MHz clock
   input reset,		// 1 to initialize module
   input sync_serial,
   input move,
	
   input [10:0] hcount,	// horizontal index of current pixel (0..1023)
   input [9:0] 	vcount, // vertical index of current pixel (0..767)
   input hsync,		// XVGA horizontal sync signal (active low)
   input vsync,		// XVGA vertical sync signal (active low)
   input blank,		// XVGA blanking (1 means output black pixel)
   input keyboard_clock, keyboard_data,
   output phsync,	// pong game's horizontal sync
   output pvsync,	// pong game's vertical sync
   output pblank,	// pong game's blanking
	output reg have_trigger,
   output [23:0] pixel,	// pong game's pixel  // r=23:16, g=15:8, b=7:0
   output [10:0]_x, 
	output [9:0] _y, output reg show_trigger, output counting
   );

   wire [2:0] checkerboard;
	
   // REPLACE ME! The code below just generates a color checkerboard
   // using 64 pixel by 64 pixel squares.
   ///Rain bow blobs parameters
   //.x(128),.x1(224),.x2(320),.x3(416)
   parameter X = 128;
   parameter X1 = 224;
   parameter X2 = 320;
   parameter X3 = 416;
   ////hit blobs
   wire [10:0] x;
   wire [9:0] y;
	reg [10:0] hit_x,_hit_x;
	reg [9:0]  hit_y, _hit_y;
	
	wire trigger, clear, ready, increase_score,_clear;
   wire [23:0] h_pixel;
   assign _x=hit_x;
	assign _y = hit_y;
	parameter TRIGGERING = 12_000_000;
	reg [26:0] trig_count;
	//reg have_trigger;
   read_ir_data receiver(.reset(reset), .clk(clk), .serial(~sync_serial),.ready(ready),.x(x), .y(y), .trigger(trigger),.clear(clear));
	always @(posedge clk) begin
	  hit_x = (ready)?x:hit_x;
	  hit_y = (ready)?y:hit_y;
	  if (ready) begin
	    if (!trigger) show_trigger <= 1;
		 have_trigger<=(trig_count>=TRIGGERING)?0:((trigger)?1:((clear)?0:0));
		 
		 
	  end
	  trig_count<=(have_trigger)?trig_count+1:0;
	  _hit_x = (ready)?x:_hit_x;
	  _hit_y = (ready)?y:_hit_y;
	  //have_trigger<=trigger;
	end 
	assign _clear = clear;
   ///
   incident_blob bullet_blobs(.x(hit_x),.y(hit_y),.hcount(hcount),.vcount(vcount),.clk(vclock),.clear(clear),
	                           .trigger(trigger),.pixel(h_pixel), .see_counting(counting), .increase_score(increase_score));
   ///////SCORE DISPLAY AREA
  wire [17:0] score_text;
  wire [23:0] score_pixel, key_pixel, text_pixel;
  wire [6:0] score;
  wire [9:0] cumm_score;
  wire [59:0] name_text;
  reg [59:0] input_text;
  wire backspace, kbd_start, enter;
  reg store_kbd_ready, store_bkspc, store_enter;
  assign score_pixel = text_pixel|key_pixel;

   multiple_text disp_score(.text(score_text), .x(466), .hcount(hcount), .y(730), .vcount(vcount),
		               .clk(vclock), .pixel(text_pixel));
   multiple_text disp_name(.text(input_text), .x(400), .y(660), .hcount(hcount), .vcount(vcount),
                           .clk(vclock), .pixel(key_pixel));

   score scr(.x(_hit_x), .center_x(512), .y(_hit_y), .center_y(384), .clk(vclock), 
		     .trigger(increase_score), .clear(_clear), .score(score), .score_text(score_text), 
		     .cumm_sc(cumm_score));

  keyboard kbd(.clk(clk), .reset(reset), .kbd_clk(keyboard_clock), .data(keyboard_data),
               .kbd_start(kbd_start), .name(name_text), .backspace(backspace), .enter(enter)); 

  reg [9:0] vertical_pose=0;
  always @(posedge vclock) begin
    if(hcount==1023&& vcount==767) begin
			
		store_kbd_ready <= kbd_start; store_bkspc <= backspace;
		store_enter <= enter;

		// update text on text input, backspace or enter
		if ((backspace != store_bkspc) || (kbd_start != store_kbd_ready)
			  || (enter != store_enter)) begin
		  input_text <= name_text;
		end

      vertical_pose<=(vertical_pose<767)?vertical_pose+2:0;
    
    end 
  end 
  wire [23:0] moving_pixel;
  leaf lf(.clk(vclock), .x(180),.hcount(hcount), .y(vertical_pose),.vcount(vcount), 
      .pixel(moving_pixel));
	/////END OF DISPLAY SCORE AREA

   /////make the circles move
   wire [23:0] xpixel;
   reg [10:0] x_0, x_1, x_2, x_3;
   reg [6:0] add_pose;
   reg right;
   reg increase;
   always @(posedge clk) begin
      if (move||(hcount==1023&&vcount==767)) begin
         add_pose<=(add_pose<=50|increase)?add_pose+1:((add_pose>=0)?add_pose-1:0);
         increase<=(add_pose==49|add_pose==49)?~increase:increase;
         right<=(add_pose==49)?!increase:increase;
         x_0<=(right)?(x_0+add_pose):(x_0-add_pose);
         x_1<=(right)?(x_1+add_pose):(x_1-add_pose);
         x_2<=(right)?(x_2+add_pose):(x_2-add_pose);
         x_3<=(right)?(x_3+add_pose):(x_3-add_pose);
     end
     else begin
       add_pose<=0;
         increase<=1;
         right<=1;
         x_0<=X;
         x_1<=X1;
         x_2<=X2;
         x_3<=X3;
     end 
   end 
////END
   circles crcls(.clk(vclock), .x(x_0),.x1(x_1),.x2(x_2),.x3(x_3), .hcount(hcount), .y(0),.y1(96),.y2(192),.y3(288), .vcount(vcount), .pixel(xpixel));
   assign phsync = hsync;
   assign pvsync = vsync;
   assign pblank = blank;
   assign checkerboard = hcount[8:6] + vcount[8:6];
   
	
	/////SOUND TRIGGER SETUP
//	reg [1:0] trig_state;
//	reg snd_trigger;
//	always @(posedge clk) begin
//	   case(trig_state)
//		  
//		endcase
//	end 
	/////////END SOUND TRIGGER SETUP
	//wire [10:0] cx;
	 //wire [9:0] cy;
	 //center_calc cenc(.clk(clk),.hcount(hcount), .vcount(vcount), .pixel(black_white), .cx(cx),.cy(cy));
	 wire [23:0] b_pixel;
	 blob bl1(.x(64),.hcount(hcount), .y(64),.vcount(hcount), .pixel(b_pixel));
   // here we use three bits from hcount and vcount to generate the \
   // checkerboard
   wire [23:0] disp_pixel;
   assign disp_pixel = (h_pixel>1)?{xpixel[23:16]>>1+h_pixel[23:16]>>1, xpixel[15:8]>>1+h_pixel[15:8]>>1,xpixel[7:0]>>1+h_pixel[7:0]>>1}:xpixel;//{{8{checkerboard[2]}}, {8{checkerboard[1]}}, {8{checkerboard[0]}}} ;
   assign pixel = (moving_pixel[23:16]>200)?moving_pixel:(score_pixel>3)?{disp_pixel[23:16]>>1+score_pixel[23:16]>>1, disp_pixel[15:8]>>1+score_pixel[15:8]>>1,disp_pixel[7:0]>>1+score_pixel[7:0]>>1}:disp_pixel;
     
endmodule

module blob
   #(parameter WIDTH = 64,            // default width: 64 pixels
               HEIGHT = 64,           // default height: 64 pixels
               COLOR = 24'hFF_FF_FF)  // default color: white
   (input [10:0] x,hcount,
    input [9:0] y,vcount,
    output reg [23:0] pixel);

   always @ * begin
      if ((hcount >= x && hcount < (x+WIDTH)) && (vcount >= y && vcount < (y+HEIGHT)))
	pixel = COLOR;
      else pixel = 0;
   end
endmodule
